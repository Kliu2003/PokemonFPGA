//module pkm_tb;
//	PokemonFPGA pkm(.*);
//	logic 
//endmodule 